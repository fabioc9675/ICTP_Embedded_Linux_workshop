----------------------------------------------------------------------------------
-- Generador de medio círculo (semicircular wave)
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity biexponential is
    Port ( 
            clk        : in  STD_LOGIC;
            rst        : in  STD_LOGIC;
            semi_out   : out STD_LOGIC_VECTOR (15 downto 0)
         );
end biexponential;

architecture Behavioral of biexponential is

    type biexponential_table is array(0 to 255) of integer range 0 to 65535;
    constant bi_exp_table : biexponential_table := (
        0, 0, 0, 0, 0, 0, 0, 0,
        0, 0, 0, 0, 0, 0, 0, 0,
        0, 0, 0, 0, 0, 0, 0, 0,
        0, 3179, 28977, 45374, 55460, 61320, 64362, 65535,
        65479, 64627, 63266, 61593, 59738, 57788, 55800, 53812,
        51850, 49928, 48057, 46242, 44486, 42790, 41154, 39579,
        38061, 36601, 35195, 33843, 32543, 31292, 30089, 28932,
        27820, 26750, 25721, 24732, 23781, 22867, 21987, 21142,
        20329, 19547, 18795, 18072, 17377, 16709, 16067, 15449,
        14855, 14283, 13734, 13206, 12698, 12210, 11740, 11289,
        10855, 10437, 10036, 9650, 9279, 8922, 8579, 8249,
        7932, 7627, 7333, 7051, 6780, 6519, 6269, 6028,
        5796, 5573, 5359, 5153, 4954, 4764, 4581, 4404,
        4235, 4072, 3916, 3765, 3620, 3481, 3347, 3218,
        3095, 2976, 2861, 2751, 2645, 2544, 2446, 2352,
        2261, 2174, 2091, 2010, 1933, 1859, 1787, 1718,
        1652, 1589, 1528, 1469, 1413, 1358, 1306, 1256,
        1207, 1161, 1116, 1073, 1032, 992, 954, 918,
        882, 848, 816, 784, 754, 725, 697, 671,
        645, 620, 596, 573, 551, 530, 510, 490,
        471, 453, 436, 419, 403, 387, 372, 358,
        344, 331, 318, 306, 294, 283, 272, 262,
        252, 242, 233, 224, 215, 207, 199, 191,
        184, 177, 170, 163, 157, 151, 145, 140,
        134, 129, 124, 119, 115, 110, 106, 102,
        98, 94, 91, 87, 84, 81, 78, 75,
        72, 69, 66, 64, 61, 59, 57, 55,
        52, 50, 48, 47, 45, 43, 41, 40,
        38, 37, 35, 34, 33, 31, 30, 29,
        28, 27, 26, 25, 24, 23, 22, 21,
        20, 20, 19, 18, 17, 17, 16, 16,
        15, 14, 14, 13, 13, 12, 12, 11
    );

    signal idx  : integer range 0 to 255 := 0;
    signal val  : integer range 0 to 65535 := 0;

begin
    process(clk, rst)
    begin
        if rst = '1' then
            idx <= 0;
            val <= bi_exp_table(0);
        elsif rising_edge(clk) then
            val <= bi_exp_table(idx);
            semi_out <= conv_std_logic_vector(val, 16);

            if idx = 255 then
                idx <= 0;
            else
                idx <= idx + 1;
            end if;
        end if;
    end process;
end Behavioral;