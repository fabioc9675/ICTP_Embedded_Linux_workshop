----------------------------------------------------------------------------------
-- Generador de medio círculo (semicircular wave)
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity semicircle_wave_gen is
    Port ( 
            clk        : in  STD_LOGIC;
            rst        : in  STD_LOGIC;
            semi_out   : out STD_LOGIC_VECTOR (15 downto 0)
         );
end semicircle_wave_gen;

architecture Behavioral of semicircle_wave_gen is

    type semicircle_table is array(0 to 255) of integer range 0 to 65535;
    constant semi_table : semicircle_table := (
        0, 8192, 11562, 14133, 16287, 18173, 19867, 21416,
        22849, 24186, 25442, 26629, 27756, 28830, 29857, 30840,
        31785, 32695, 33572, 34419, 35238, 36032, 36801, 37547,
        38272, 38976, 39662, 40329, 40979, 41612, 42230, 42832,
        43420, 43995, 44556, 45104, 45639, 46163, 46675, 47176,
        47667, 48147, 48616, 49076, 49526, 49967, 50399, 50821,
        51236, 51641, 52039, 52428, 52810, 53184, 53550, 53909,
        54261, 54606, 54943, 55274, 55598, 55916, 56226, 56531,
        56829, 57122, 57408, 57688, 57962, 58230, 58493, 58750,
        59001, 59247, 59487, 59722, 59951, 60176, 60395, 60609,
        60818, 61022, 61220, 61414, 61603, 61787, 61967, 62141,
        62311, 62476, 62637, 62793, 62944, 63091, 63233, 63371,
        63504, 63633, 63757, 63877, 63993, 64104, 64211, 64314,
        64413, 64507, 64597, 64683, 64764, 64842, 64915, 64984,
        65049, 65110, 65167, 65220, 65268, 65313, 65353, 65390,
        65422, 65450, 65475, 65495, 65511, 65523, 65531, 65535,
        65535, 65531, 65523, 65511, 65495, 65475, 65450, 65422,
        65390, 65353, 65313, 65268, 65220, 65167, 65110, 65049,
        64984, 64915, 64842, 64764, 64683, 64597, 64507, 64413,
        64314, 64211, 64104, 63993, 63877, 63757, 63633, 63504,
        63371, 63233, 63091, 62944, 62793, 62637, 62476, 62311,
        62141, 61967, 61787, 61603, 61414, 61220, 61022, 60818,
        60609, 60395, 60176, 59951, 59722, 59487, 59247, 59001,
        58750, 58493, 58230, 57962, 57688, 57408, 57122, 56829,
        56531, 56226, 55916, 55598, 55274, 54943, 54606, 54261,
        53909, 53550, 53184, 52810, 52428, 52039, 51641, 51236,
        50821, 50399, 49967, 49526, 49076, 48616, 48147, 47667,
        47176, 46675, 46163, 45639, 45104, 44556, 43995, 43420,
        42832, 42230, 41612, 40979, 40329, 39662, 38976, 38272,
        37547, 36801, 36032, 35238, 34419, 33572, 32695, 31785,
        30840, 29857, 28830, 27756, 26629, 25442, 24186, 22849,
        21416, 19867, 18173, 16287, 14133, 11562, 8192, 0
    );

    signal idx  : integer range 0 to 255 := 0;
    signal val  : integer range 0 to 65535 := 0;

begin
    process(clk, rst)
    begin
        if rst = '1' then
            idx <= 0;
            val <= semi_table(0);
        elsif rising_edge(clk) then
            val <= semi_table(idx);
            semi_out <= conv_std_logic_vector(val, 16);

            if idx = 255 then
                idx <= 0;
            else
                idx <= idx + 1;
            end if;
        end if;
    end process;
end Behavioral;